* dual rc ladder
R1 int in 10k
V1 in 0 dc 0 PULSE (0 5 1u 1u 1u 1 1)
R2 out int 1k
C1 int 0 1u
C2 out 0 100n
* .option trtol=1 klu method=gear reltol=1m
* .option sparse
.tran 50u 200u 0 0.1u
.save v(in) v(int) v(out)
.end